**************************************************
* ����ģ���·����������ϵͳ������·��             *
**************************************************
* �����������¿������ܽ�                       *
**************************************************
* �������� ��ѧ�����硡2020                      *
**************************************************

.SUBCKT CS_AMP GNDA VDDA vin vout Vbias

* with current-source load
MM1 vout vin	 GNDA GNDA n18	W=10u	L=180n	M=1
MM2 vout Vbias VDDA VDDA p18	W=60u	L=1u	M=1

.ENDS