﻿**************************************************
* 　　模拟电路基础——从系统级到电路级             *
**************************************************
* 　　　　　陈抗生　周金芳                       *
**************************************************
* 　　　　 科学出版社　2020                      *
**************************************************          

.title book_6.5


.param W1=5u
M1 2 1 0 0 n18 W=W1 L=180n m=1
VVDS 2 0 DC 1.8V
VVGS 1 0 DC 0.75V

.op
.dc VVDS 0 1.8 0.1 W1 5u 25u 5u

.print gm=lx7(M1) gds=lx8(M1) cgs=par('-lx20(M1)') cgd=par('-lx19(M1)') 

.probe v(2) v(1) i(M1)

.temp 27
.option post accurate probe
.lib '..\models\ms018.lib' tt

.end