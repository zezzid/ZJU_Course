﻿**************************************************
* 　　模拟电路基础——从系统级到电路级             *
**************************************************
* 　　　　　陈抗生　周金芳                       *
**************************************************
* 　　　　 科学出版社　2020                      *
**************************************************          

.title NMOS_DC

VVDS net2 0 DC 1.8V
VVGS net1 0 DC 0.75V
MNM0 net2 net1 0 0 n18 W=5u L=180n m=1

.op                                 * 打印直流工作点
.dc VVDS 0 1.8 0.1 VVGS 0 1.8 0.3   * 直流仿真，设置扫描变量，
                                    * 范围0-1.8V，步长分别为0.1V和0.3V
.probe v(net2) v(net1) i(MNM0)

.temp 27
.option post accurate probe
.lib '..\models\ms018.lib' tt

.end